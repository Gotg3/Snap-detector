library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

	entity snap_dec_tx_mic_tb is
	end snap_dec_tx_mic_tb;
	
	
	architecture dut of snap_dec_tx_mic_tb is
	
	
	component snap_dec_mic
	port(
		pdm: in std_logic; -- ingresso pdm 
		--pdm_in_dx: in std_logic; -- ingresso pdm canale dx
		--decision: out std_logic_vector(7 downto 0);
		clk: in std_logic;
		rst: in std_logic;
		ack: in std_logic; --ack che arriva alla uart
		TX: out std_logic -- uscita seriale della UART
		);
	end component;
	
	--signal pdm: std_logic;
	--signal pdm_dx_sig: std_logic;
	signal clk_sig: std_logic:='0';
	signal rst_sig: std_logic;
	signal ack_sig: std_logic;  -- messo a uno così trasmette con continuità, è una prova..
	signal TX_sig: std_logic;
	signal clk_demux: std_logic:='0';
	signal vect1_PDM : std_logic_vector(0 to 3374):="010101101010101010101010101010101010101010101010101010101010100101010101010101010010101010101010010101010101010100101010101010101010101010101010101010101010101011010101010101010110101010101010110101010101101010101011010101011010101011010101011010101011010101101010110101011010101101010101101010110101011010101011010101101010101101010101011010101010110101010101011010101010101011010101010101010101011010101010101010101010101010101010101010101010100101010101010101001010101010100101010100101010100101010100101010100101010101001010101001010101010100101010101010101010101010101010101010101010110101010101101010110101011010110101101011011010110110110110110110110110111011011101101110111011011101110111011101110111011110111011101110111011101110111011101101110111011011101101110110110110110110110110110110110110110101101011011010101101011010101101010101010110101010101010101010101010101010100101010101010101010010101010101010010101010101010010101010101010101001010101010101010101010101010101010101010101010101010101010110101010101101010101101010110101011010101101010110101011010101101010110101010110101010110101010110101010110101010110101010110101011010101011010101101010110101011010101101010101101010110101011010101011010101011010101010110101010101011010101010101010101010101010101010101010100101010100101010100101001010100101001010010010100100101001001001001001001001001001001001001000100100010010001000100010001000100010001000010001000010000100010000100001000001000010000100001000010001000010000100010000100010001000100010001000100010001001000100010010010001001000100100100100010010010010010010010010010010010010100100100101001001010010010100101001010100101010010101001010101010100101010101010101010101010101010101011010101010101101010110101011010101101011010110101101011010110110101101101101011011011011011011011011011011011011011011101101101110110110111011011101101110111011011101101110111011011101110110111011101101110110111011011101101101110110111011011011101101101110110110110111011011011011101101101101101101101101110110101101101101101101101011011010110110101101011010110101101011010101101010110101011010101010110101010101101010101010101010101010101010101010101010101001010101010010101010010101001010010101001010010100101010010100101001010010100101001010010100101001010010100101001010010100101001010100101001010010100101010010100101010010100101010010100101010010100101010010100101001010100101001010010100101001010010100101001010010010100101001001010010100100101001001010010010100100100101001001001001001001010010010010010010010010010010010010010010010010010010010010010010100100100100101001001010010100101001010010101001010100101010101001010101010101010101010101010101010101010101010101011010101010101101010101011010101011010101011010101011010101011010101101010101101010101101010110101011010101011010101011010101101010101101010101011010101011010101010101101010101010110101010101010110101010101010110101010101010110101010101011010101010110101010110101011010101101010110101101011010110101101011010110110101101101011011010110110110101101101011011011010110110110101101101011011011010110110101101101011010110110101101011010110101101011010110101101011010101101010110101011010101011010101011010101010101011010101010101010101010101010101010101010101010010101010101010101001010101010101001010101010100101010101010010101010101001010101010010101010100101010101001010101001010101010010";
	
	signal vect1_PDM_noise: std_logic_vector(0 to 3374):="101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101";
	signal PDM_sig: std_logic;
signal pdm_dx_sig: std_logic;
signal pdm_sx_sig: std_logic;
		
	
	begin
	
	sn_tx: component snap_dec_mic
	port map(
	pdm=>PDM_sig,
	clk=>clk_sig,
	rst=>rst_sig,
	ack=>ack_sig,
	TX=>TX_sig
	);
	
	
	clk_sig<= not(clk_sig) after 20 ns; --periodo di 25Mhz (semiperiodo di 20 ns)
	clk_demux<=not(clk_demux) after 520 ns; -- clock a 4 MHz per ddr
	
	mux_cod: process(clk_demux,pdm_dx_sig,pdm_sx_sig) --codifica il pdm
	begin					 
		if (clk_demux='1') then	
			PDM_sig<=pdm_dx_sig;
		else
			PDM_sig<=pdm_sx_sig;
		end if;
	end process;
	

	
	
	
	stimuli: process
	
	begin 
	ack_sig<='1';
	rst_sig <= '1','0' after 40 ns;
	
		for k in 0 to 3374 loop 
		
		pdm_dx_sig <=vect1_PDM_noise(k) ; 
       		 pdm_sx_sig <=vect1_PDM(k) ;
		wait for 520 ns;
		end loop ;
	
        for k in 0 to 3374 loop 
        pdm_dx_sig <=vect1_PDM_noise(k) ; 
        pdm_sx_sig <=vect1_PDM(k) ; 
		
        wait for 520 ns;
        end loop ;
		
		for k in 0 to 3374 loop  
        pdm_dx_sig <=vect1_PDM_noise(k) ; 
        pdm_sx_sig <=vect1_PDM_noise(k) ; 
        wait for 520 ns;
        end loop ;


--------
	





    pdm_dx_sig <='0';
	pdm_sx_sig <='0';


	
	wait;

	end process;

end architecture;
	
	